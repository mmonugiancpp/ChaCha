/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_mmonugiancpp (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  assign uio_oe = 8'b11111000;

  ChaChaEncryption mybaby(
                clk,
                ~rst_n,
                0,
                0,
                0,
                0,
                0,
                0,
                0,
                0,
                0,
                0,
                0,
                0,
                uio_in[0],
                ui_in,
                uio_in[1],
                uio_out[3],
                uo_out,
                uio_out[4],
                uio_in[2]
  );
  // All output pins must be assigned. If not used, assign to 0.
  assign uio_out[7:5] = 3'b000;
  assign uio_out[2:0] = 3'b000;

  // List all unused inputs to prevent warnings
    wire _unused = &{uio_in[7:3], 1'b0};

endmodule


